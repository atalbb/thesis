`timescale 10ns / 1ps

module mixcolumn(a,mcl,decrypt);
input [127:0] a;
input decrypt;
output [127:0] mcl;

assign mcl = (decrypt==0)?mixcolumns(a):inv_mixcolumns(a);

//wire [7 : 0] mul2 [0 : 255];
//wire [7 : 0] mul3 [0 : 255];
//wire [7 : 0] mul9 [0 : 255];
//wire [7 : 0] mul11 [0 : 255];
//wire [7 : 0] mul13 [0 : 255];
//wire [7 : 0] mul14 [0 : 255];

//assign mul2[8'h00] = 8'h00;
//assign mul2[8'h01] = 8'h02;
//assign mul2[8'h02] = 8'h04;
//assign mul2[8'h03] = 8'h06;
//assign mul2[8'h04] = 8'h08;
//assign mul2[8'h05] = 8'h0a;
//assign mul2[8'h06] = 8'h0c;
//assign mul2[8'h07] = 8'h0e;
//assign mul2[8'h08] = 8'h10;
//assign mul2[8'h09] = 8'h12;
//assign mul2[8'h0a] = 8'h14;
//assign mul2[8'h0b] = 8'h16;
//assign mul2[8'h0c] = 8'h18;
//assign mul2[8'h0d] = 8'h1a;
//assign mul2[8'h0e] = 8'h1c;
//assign mul2[8'h0f] = 8'h1e;
//assign mul2[8'h10] = 8'h20;
//assign mul2[8'h11] = 8'h22;
//assign mul2[8'h12] = 8'h24;
//assign mul2[8'h13] = 8'h26;
//assign mul2[8'h14] = 8'h28;
//assign mul2[8'h15] = 8'h2a;
//assign mul2[8'h16] = 8'h2c;
//assign mul2[8'h17] = 8'h2e;
//assign mul2[8'h18] = 8'h30;
//assign mul2[8'h19] = 8'h32;
//assign mul2[8'h1a] = 8'h34;
//assign mul2[8'h1b] = 8'h36;
//assign mul2[8'h1c] = 8'h38;
//assign mul2[8'h1d] = 8'h3a;
//assign mul2[8'h1e] = 8'h3c;
//assign mul2[8'h1f] = 8'h3e;
//assign mul2[8'h20] = 8'h40;
//assign mul2[8'h21] = 8'h42;
//assign mul2[8'h22] = 8'h44;
//assign mul2[8'h23] = 8'h46;
//assign mul2[8'h24] = 8'h48;
//assign mul2[8'h25] = 8'h4a;
//assign mul2[8'h26] = 8'h4c;
//assign mul2[8'h27] = 8'h4e;
//assign mul2[8'h28] = 8'h50;
//assign mul2[8'h29] = 8'h52;
//assign mul2[8'h2a] = 8'h54;
//assign mul2[8'h2b] = 8'h56;
//assign mul2[8'h2c] = 8'h58;
//assign mul2[8'h2d] = 8'h5a;
//assign mul2[8'h2e] = 8'h5c;
//assign mul2[8'h2f] = 8'h5e;
//assign mul2[8'h30] = 8'h60;
//assign mul2[8'h31] = 8'h62;
//assign mul2[8'h32] = 8'h64;
//assign mul2[8'h33] = 8'h66;
//assign mul2[8'h34] = 8'h68;
//assign mul2[8'h35] = 8'h6a;
//assign mul2[8'h36] = 8'h6c;
//assign mul2[8'h37] = 8'h6e;
//assign mul2[8'h38] = 8'h70;
//assign mul2[8'h39] = 8'h72;
//assign mul2[8'h3a] = 8'h74;
//assign mul2[8'h3b] = 8'h76;
//assign mul2[8'h3c] = 8'h78;
//assign mul2[8'h3d] = 8'h7a;
//assign mul2[8'h3e] = 8'h7c;
//assign mul2[8'h3f] = 8'h7e;
//assign mul2[8'h40] = 8'h80;
//assign mul2[8'h41] = 8'h82;
//assign mul2[8'h42] = 8'h84;
//assign mul2[8'h43] = 8'h86;
//assign mul2[8'h44] = 8'h88;
//assign mul2[8'h45] = 8'h8a;
//assign mul2[8'h46] = 8'h8c;
//assign mul2[8'h47] = 8'h8e;
//assign mul2[8'h48] = 8'h90;
//assign mul2[8'h49] = 8'h92;
//assign mul2[8'h4a] = 8'h94;
//assign mul2[8'h4b] = 8'h96;
//assign mul2[8'h4c] = 8'h98;
//assign mul2[8'h4d] = 8'h9a;
//assign mul2[8'h4e] = 8'h9c;
//assign mul2[8'h4f] = 8'h9e;
//assign mul2[8'h50] = 8'ha0;
//assign mul2[8'h51] = 8'ha2;
//assign mul2[8'h52] = 8'ha4;
//assign mul2[8'h53] = 8'ha6;
//assign mul2[8'h54] = 8'ha8;
//assign mul2[8'h55] = 8'haa;
//assign mul2[8'h56] = 8'hac;
//assign mul2[8'h57] = 8'hae;
//assign mul2[8'h58] = 8'hb0;
//assign mul2[8'h59] = 8'hb2;
//assign mul2[8'h5a] = 8'hb4;
//assign mul2[8'h5b] = 8'hb6;
//assign mul2[8'h5c] = 8'hb8;
//assign mul2[8'h5d] = 8'hba;
//assign mul2[8'h5e] = 8'hbc;
//assign mul2[8'h5f] = 8'hbe;
//assign mul2[8'h60] = 8'hc0;
//assign mul2[8'h61] = 8'hc2;
//assign mul2[8'h62] = 8'hc4;
//assign mul2[8'h63] = 8'hc6;
//assign mul2[8'h64] = 8'hc8;
//assign mul2[8'h65] = 8'hca;
//assign mul2[8'h66] = 8'hcc;
//assign mul2[8'h67] = 8'hce;
//assign mul2[8'h68] = 8'hd0;
//assign mul2[8'h69] = 8'hd2;
//assign mul2[8'h6a] = 8'hd4;
//assign mul2[8'h6b] = 8'hd6;
//assign mul2[8'h6c] = 8'hd8;
//assign mul2[8'h6d] = 8'hda;
//assign mul2[8'h6e] = 8'hdc;
//assign mul2[8'h6f] = 8'hde;
//assign mul2[8'h70] = 8'he0;
//assign mul2[8'h71] = 8'he2;
//assign mul2[8'h72] = 8'he4;
//assign mul2[8'h73] = 8'he6;
//assign mul2[8'h74] = 8'he8;
//assign mul2[8'h75] = 8'hea;
//assign mul2[8'h76] = 8'hec;
//assign mul2[8'h77] = 8'hee;
//assign mul2[8'h78] = 8'hf0;
//assign mul2[8'h79] = 8'hf2;
//assign mul2[8'h7a] = 8'hf4;
//assign mul2[8'h7b] = 8'hf6;
//assign mul2[8'h7c] = 8'hf8;
//assign mul2[8'h7d] = 8'hfa;
//assign mul2[8'h7e] = 8'hfc;
//assign mul2[8'h7f] = 8'hfe;
//assign mul2[8'h80] = 8'h1b;
//assign mul2[8'h81] = 8'h19;
//assign mul2[8'h82] = 8'h1f;
//assign mul2[8'h83] = 8'h1d;
//assign mul2[8'h84] = 8'h13;
//assign mul2[8'h85] = 8'h11;
//assign mul2[8'h86] = 8'h17;
//assign mul2[8'h87] = 8'h15;
//assign mul2[8'h88] = 8'h0b;
//assign mul2[8'h89] = 8'h09;
//assign mul2[8'h8a] = 8'h0f;
//assign mul2[8'h8b] = 8'h0d;
//assign mul2[8'h8c] = 8'h03;
//assign mul2[8'h8d] = 8'h01;
//assign mul2[8'h8e] = 8'h07;
//assign mul2[8'h8f] = 8'h05;
//assign mul2[8'h90] = 8'h3b;
//assign mul2[8'h91] = 8'h39;
//assign mul2[8'h92] = 8'h3f;
//assign mul2[8'h93] = 8'h3d;
//assign mul2[8'h94] = 8'h33;
//assign mul2[8'h95] = 8'h31;
//assign mul2[8'h96] = 8'h37;
//assign mul2[8'h97] = 8'h35;
//assign mul2[8'h98] = 8'h2b;
//assign mul2[8'h99] = 8'h29;
//assign mul2[8'h9a] = 8'h2f;
//assign mul2[8'h9b] = 8'h2d;
//assign mul2[8'h9c] = 8'h23;
//assign mul2[8'h9d] = 8'h21;
//assign mul2[8'h9e] = 8'h27;
//assign mul2[8'h9f] = 8'h25;
//assign mul2[8'ha0] = 8'h5b;
//assign mul2[8'ha1] = 8'h59;
//assign mul2[8'ha2] = 8'h5f;
//assign mul2[8'ha3] = 8'h5d;
//assign mul2[8'ha4] = 8'h53;
//assign mul2[8'ha5] = 8'h51;
//assign mul2[8'ha6] = 8'h57;
//assign mul2[8'ha7] = 8'h55;
//assign mul2[8'ha8] = 8'h4b;
//assign mul2[8'ha9] = 8'h49;
//assign mul2[8'haa] = 8'h4f;
//assign mul2[8'hab] = 8'h4d;
//assign mul2[8'hac] = 8'h43;
//assign mul2[8'had] = 8'h41;
//assign mul2[8'hae] = 8'h47;
//assign mul2[8'haf] = 8'h45;
//assign mul2[8'hb0] = 8'h7b;
//assign mul2[8'hb1] = 8'h79;
//assign mul2[8'hb2] = 8'h7f;
//assign mul2[8'hb3] = 8'h7d;
//assign mul2[8'hb4] = 8'h73;
//assign mul2[8'hb5] = 8'h71;
//assign mul2[8'hb6] = 8'h77;
//assign mul2[8'hb7] = 8'h75;
//assign mul2[8'hb8] = 8'h6b;
//assign mul2[8'hb9] = 8'h69;
//assign mul2[8'hba] = 8'h6f;
//assign mul2[8'hbb] = 8'h6d;
//assign mul2[8'hbc] = 8'h63;
//assign mul2[8'hbd] = 8'h61;
//assign mul2[8'hbe] = 8'h67;
//assign mul2[8'hbf] = 8'h65;
//assign mul2[8'hc0] = 8'h9b;
//assign mul2[8'hc1] = 8'h99;
//assign mul2[8'hc2] = 8'h9f;
//assign mul2[8'hc3] = 8'h9d;
//assign mul2[8'hc4] = 8'h93;
//assign mul2[8'hc5] = 8'h91;
//assign mul2[8'hc6] = 8'h97;
//assign mul2[8'hc7] = 8'h95;
//assign mul2[8'hc8] = 8'h8b;
//assign mul2[8'hc9] = 8'h89;
//assign mul2[8'hca] = 8'h8f;
//assign mul2[8'hcb] = 8'h8d;
//assign mul2[8'hcc] = 8'h83;
//assign mul2[8'hcd] = 8'h81;
//assign mul2[8'hce] = 8'h87;
//assign mul2[8'hcf] = 8'h85;
//assign mul2[8'hd0] = 8'hbb;
//assign mul2[8'hd1] = 8'hb9;
//assign mul2[8'hd2] = 8'hbf;
//assign mul2[8'hd3] = 8'hbd;
//assign mul2[8'hd4] = 8'hb3;
//assign mul2[8'hd5] = 8'hb1;
//assign mul2[8'hd6] = 8'hb7;
//assign mul2[8'hd7] = 8'hb5;
//assign mul2[8'hd8] = 8'hab;
//assign mul2[8'hd9] = 8'ha9;
//assign mul2[8'hda] = 8'haf;
//assign mul2[8'hdb] = 8'had;
//assign mul2[8'hdc] = 8'ha3;
//assign mul2[8'hdd] = 8'ha1;
//assign mul2[8'hde] = 8'ha7;
//assign mul2[8'hdf] = 8'ha5;
//assign mul2[8'he0] = 8'hdb;
//assign mul2[8'he1] = 8'hd9;
//assign mul2[8'he2] = 8'hdf;
//assign mul2[8'he3] = 8'hdd;
//assign mul2[8'he4] = 8'hd3;
//assign mul2[8'he5] = 8'hd1;
//assign mul2[8'he6] = 8'hd7;
//assign mul2[8'he7] = 8'hd5;
//assign mul2[8'he8] = 8'hcb;
//assign mul2[8'he9] = 8'hc9;
//assign mul2[8'hea] = 8'hcf;
//assign mul2[8'heb] = 8'hcd;
//assign mul2[8'hec] = 8'hc3;
//assign mul2[8'hed] = 8'hc1;
//assign mul2[8'hee] = 8'hc7;
//assign mul2[8'hef] = 8'hc5;
//assign mul2[8'hf0] = 8'hfb;
//assign mul2[8'hf1] = 8'hf9;
//assign mul2[8'hf2] = 8'hff;
//assign mul2[8'hf3] = 8'hfd;
//assign mul2[8'hf4] = 8'hf3;
//assign mul2[8'hf5] = 8'hf1;
//assign mul2[8'hf6] = 8'hf7;
//assign mul2[8'hf7] = 8'hf5;
//assign mul2[8'hf8] = 8'heb;
//assign mul2[8'hf9] = 8'he9;
//assign mul2[8'hfa] = 8'hef;
//assign mul2[8'hfb] = 8'hed;
//assign mul2[8'hfc] = 8'he3;
//assign mul2[8'hfd] = 8'he1;
//assign mul2[8'hfe] = 8'he7;
//assign mul2[8'hff] = 8'he5;

//assign mul3[8'h00] = 8'h00;
//assign mul3[8'h01] = 8'h03;
//assign mul3[8'h02] = 8'h06;
//assign mul3[8'h03] = 8'h05;
//assign mul3[8'h04] = 8'h0c;
//assign mul3[8'h05] = 8'h0f;
//assign mul3[8'h06] = 8'h0a;
//assign mul3[8'h07] = 8'h09;
//assign mul3[8'h08] = 8'h18;
//assign mul3[8'h09] = 8'h1b;
//assign mul3[8'h0a] = 8'h1e;
//assign mul3[8'h0b] = 8'h1d;
//assign mul3[8'h0c] = 8'h14;
//assign mul3[8'h0d] = 8'h17;
//assign mul3[8'h0e] = 8'h12;
//assign mul3[8'h0f] = 8'h11;
//assign mul3[8'h10] = 8'h30;
//assign mul3[8'h11] = 8'h33;
//assign mul3[8'h12] = 8'h36;
//assign mul3[8'h13] = 8'h35;
//assign mul3[8'h14] = 8'h3c;
//assign mul3[8'h15] = 8'h3f;
//assign mul3[8'h16] = 8'h3a;
//assign mul3[8'h17] = 8'h39;
//assign mul3[8'h18] = 8'h28;
//assign mul3[8'h19] = 8'h2b;
//assign mul3[8'h1a] = 8'h2e;
//assign mul3[8'h1b] = 8'h2d;
//assign mul3[8'h1c] = 8'h24;
//assign mul3[8'h1d] = 8'h27;
//assign mul3[8'h1e] = 8'h22;
//assign mul3[8'h1f] = 8'h21;
//assign mul3[8'h20] = 8'h60;
//assign mul3[8'h21] = 8'h63;
//assign mul3[8'h22] = 8'h66;
//assign mul3[8'h23] = 8'h65;
//assign mul3[8'h24] = 8'h6c;
//assign mul3[8'h25] = 8'h6f;
//assign mul3[8'h26] = 8'h6a;
//assign mul3[8'h27] = 8'h69;
//assign mul3[8'h28] = 8'h78;
//assign mul3[8'h29] = 8'h7b;
//assign mul3[8'h2a] = 8'h7e;
//assign mul3[8'h2b] = 8'h7d;
//assign mul3[8'h2c] = 8'h74;
//assign mul3[8'h2d] = 8'h77;
//assign mul3[8'h2e] = 8'h72;
//assign mul3[8'h2f] = 8'h71;
//assign mul3[8'h30] = 8'h50;
//assign mul3[8'h31] = 8'h53;
//assign mul3[8'h32] = 8'h56;
//assign mul3[8'h33] = 8'h55;
//assign mul3[8'h34] = 8'h5c;
//assign mul3[8'h35] = 8'h5f;
//assign mul3[8'h36] = 8'h5a;
//assign mul3[8'h37] = 8'h59;
//assign mul3[8'h38] = 8'h48;
//assign mul3[8'h39] = 8'h4b;
//assign mul3[8'h3a] = 8'h4e;
//assign mul3[8'h3b] = 8'h4d;
//assign mul3[8'h3c] = 8'h44;
//assign mul3[8'h3d] = 8'h47;
//assign mul3[8'h3e] = 8'h42;
//assign mul3[8'h3f] = 8'h41;
//assign mul3[8'h40] = 8'hc0;
//assign mul3[8'h41] = 8'hc3;
//assign mul3[8'h42] = 8'hc6;
//assign mul3[8'h43] = 8'hc5;
//assign mul3[8'h44] = 8'hcc;
//assign mul3[8'h45] = 8'hcf;
//assign mul3[8'h46] = 8'hca;
//assign mul3[8'h47] = 8'hc9;
//assign mul3[8'h48] = 8'hd8;
//assign mul3[8'h49] = 8'hdb;
//assign mul3[8'h4a] = 8'hde;
//assign mul3[8'h4b] = 8'hdd;
//assign mul3[8'h4c] = 8'hd4;
//assign mul3[8'h4d] = 8'hd7;
//assign mul3[8'h4e] = 8'hd2;
//assign mul3[8'h4f] = 8'hd1;
//assign mul3[8'h50] = 8'hf0;
//assign mul3[8'h51] = 8'hf3;
//assign mul3[8'h52] = 8'hf6;
//assign mul3[8'h53] = 8'hf5;
//assign mul3[8'h54] = 8'hfc;
//assign mul3[8'h55] = 8'hff;
//assign mul3[8'h56] = 8'hfa;
//assign mul3[8'h57] = 8'hf9;
//assign mul3[8'h58] = 8'he8;
//assign mul3[8'h59] = 8'heb;
//assign mul3[8'h5a] = 8'hee;
//assign mul3[8'h5b] = 8'hed;
//assign mul3[8'h5c] = 8'he4;
//assign mul3[8'h5d] = 8'he7;
//assign mul3[8'h5e] = 8'he2;
//assign mul3[8'h5f] = 8'he1;
//assign mul3[8'h60] = 8'ha0;
//assign mul3[8'h61] = 8'ha3;
//assign mul3[8'h62] = 8'ha6;
//assign mul3[8'h63] = 8'ha5;
//assign mul3[8'h64] = 8'hac;
//assign mul3[8'h65] = 8'haf;
//assign mul3[8'h66] = 8'haa;
//assign mul3[8'h67] = 8'ha9;
//assign mul3[8'h68] = 8'hb8;
//assign mul3[8'h69] = 8'hbb;
//assign mul3[8'h6a] = 8'hbe;
//assign mul3[8'h6b] = 8'hbd;
//assign mul3[8'h6c] = 8'hb4;
//assign mul3[8'h6d] = 8'hb7;
//assign mul3[8'h6e] = 8'hb2;
//assign mul3[8'h6f] = 8'hb1;
//assign mul3[8'h70] = 8'h90;
//assign mul3[8'h71] = 8'h93;
//assign mul3[8'h72] = 8'h96;
//assign mul3[8'h73] = 8'h95;
//assign mul3[8'h74] = 8'h9c;
//assign mul3[8'h75] = 8'h9f;
//assign mul3[8'h76] = 8'h9a;
//assign mul3[8'h77] = 8'h99;
//assign mul3[8'h78] = 8'h88;
//assign mul3[8'h79] = 8'h8b;
//assign mul3[8'h7a] = 8'h8e;
//assign mul3[8'h7b] = 8'h8d;
//assign mul3[8'h7c] = 8'h84;
//assign mul3[8'h7d] = 8'h87;
//assign mul3[8'h7e] = 8'h82;
//assign mul3[8'h7f] = 8'h81;
//assign mul3[8'h80] = 8'h9b;
//assign mul3[8'h81] = 8'h98;
//assign mul3[8'h82] = 8'h9d;
//assign mul3[8'h83] = 8'h9e;
//assign mul3[8'h84] = 8'h97;
//assign mul3[8'h85] = 8'h94;
//assign mul3[8'h86] = 8'h91;
//assign mul3[8'h87] = 8'h92;
//assign mul3[8'h88] = 8'h83;
//assign mul3[8'h89] = 8'h80;
//assign mul3[8'h8a] = 8'h85;
//assign mul3[8'h8b] = 8'h86;
//assign mul3[8'h8c] = 8'h8f;
//assign mul3[8'h8d] = 8'h8c;
//assign mul3[8'h8e] = 8'h89;
//assign mul3[8'h8f] = 8'h8a;
//assign mul3[8'h90] = 8'hab;
//assign mul3[8'h91] = 8'ha8;
//assign mul3[8'h92] = 8'had;
//assign mul3[8'h93] = 8'hae;
//assign mul3[8'h94] = 8'ha7;
//assign mul3[8'h95] = 8'ha4;
//assign mul3[8'h96] = 8'ha1;
//assign mul3[8'h97] = 8'ha2;
//assign mul3[8'h98] = 8'hb3;
//assign mul3[8'h99] = 8'hb0;
//assign mul3[8'h9a] = 8'hb5;
//assign mul3[8'h9b] = 8'hb6;
//assign mul3[8'h9c] = 8'hbf;
//assign mul3[8'h9d] = 8'hbc;
//assign mul3[8'h9e] = 8'hb9;
//assign mul3[8'h9f] = 8'hba;
//assign mul3[8'ha0] = 8'hfb;
//assign mul3[8'ha1] = 8'hf8;
//assign mul3[8'ha2] = 8'hfd;
//assign mul3[8'ha3] = 8'hfe;
//assign mul3[8'ha4] = 8'hf7;
//assign mul3[8'ha5] = 8'hf4;
//assign mul3[8'ha6] = 8'hf1;
//assign mul3[8'ha7] = 8'hf2;
//assign mul3[8'ha8] = 8'he3;
//assign mul3[8'ha9] = 8'he0;
//assign mul3[8'haa] = 8'he5;
//assign mul3[8'hab] = 8'he6;
//assign mul3[8'hac] = 8'hef;
//assign mul3[8'had] = 8'hec;
//assign mul3[8'hae] = 8'he9;
//assign mul3[8'haf] = 8'hea;
//assign mul3[8'hb0] = 8'hcb;
//assign mul3[8'hb1] = 8'hc8;
//assign mul3[8'hb2] = 8'hcd;
//assign mul3[8'hb3] = 8'hce;
//assign mul3[8'hb4] = 8'hc7;
//assign mul3[8'hb5] = 8'hc4;
//assign mul3[8'hb6] = 8'hc1;
//assign mul3[8'hb7] = 8'hc2;
//assign mul3[8'hb8] = 8'hd3;
//assign mul3[8'hb9] = 8'hd0;
//assign mul3[8'hba] = 8'hd5;
//assign mul3[8'hbb] = 8'hd6;
//assign mul3[8'hbc] = 8'hdf;
//assign mul3[8'hbd] = 8'hdc;
//assign mul3[8'hbe] = 8'hd9;
//assign mul3[8'hbf] = 8'hda;
//assign mul3[8'hc0] = 8'h5b;
//assign mul3[8'hc1] = 8'h58;
//assign mul3[8'hc2] = 8'h5d;
//assign mul3[8'hc3] = 8'h5e;
//assign mul3[8'hc4] = 8'h57;
//assign mul3[8'hc5] = 8'h54;
//assign mul3[8'hc6] = 8'h51;
//assign mul3[8'hc7] = 8'h52;
//assign mul3[8'hc8] = 8'h43;
//assign mul3[8'hc9] = 8'h40;
//assign mul3[8'hca] = 8'h45;
//assign mul3[8'hcb] = 8'h46;
//assign mul3[8'hcc] = 8'h4f;
//assign mul3[8'hcd] = 8'h4c;
//assign mul3[8'hce] = 8'h49;
//assign mul3[8'hcf] = 8'h4a;
//assign mul3[8'hd0] = 8'h6b;
//assign mul3[8'hd1] = 8'h68;
//assign mul3[8'hd2] = 8'h6d;
//assign mul3[8'hd3] = 8'h6e;
//assign mul3[8'hd4] = 8'h67;
//assign mul3[8'hd5] = 8'h64;
//assign mul3[8'hd6] = 8'h61;
//assign mul3[8'hd7] = 8'h62;
//assign mul3[8'hd8] = 8'h73;
//assign mul3[8'hd9] = 8'h70;
//assign mul3[8'hda] = 8'h75;
//assign mul3[8'hdb] = 8'h76;
//assign mul3[8'hdc] = 8'h7f;
//assign mul3[8'hdd] = 8'h7c;
//assign mul3[8'hde] = 8'h79;
//assign mul3[8'hdf] = 8'h7a;
//assign mul3[8'he0] = 8'h3b;
//assign mul3[8'he1] = 8'h38;
//assign mul3[8'he2] = 8'h3d;
//assign mul3[8'he3] = 8'h3e;
//assign mul3[8'he4] = 8'h37;
//assign mul3[8'he5] = 8'h34;
//assign mul3[8'he6] = 8'h31;
//assign mul3[8'he7] = 8'h32;
//assign mul3[8'he8] = 8'h23;
//assign mul3[8'he9] = 8'h20;
//assign mul3[8'hea] = 8'h25;
//assign mul3[8'heb] = 8'h26;
//assign mul3[8'hec] = 8'h2f;
//assign mul3[8'hed] = 8'h2c;
//assign mul3[8'hee] = 8'h29;
//assign mul3[8'hef] = 8'h2a;
//assign mul3[8'hf0] = 8'h0b;
//assign mul3[8'hf1] = 8'h08;
//assign mul3[8'hf2] = 8'h0d;
//assign mul3[8'hf3] = 8'h0e;
//assign mul3[8'hf4] = 8'h07;
//assign mul3[8'hf5] = 8'h04;
//assign mul3[8'hf6] = 8'h01;
//assign mul3[8'hf7] = 8'h02;
//assign mul3[8'hf8] = 8'h13;
//assign mul3[8'hf9] = 8'h10;
//assign mul3[8'hfa] = 8'h15;
//assign mul3[8'hfb] = 8'h16;
//assign mul3[8'hfc] = 8'h1f;
//assign mul3[8'hfd] = 8'h1c;
//assign mul3[8'hfe] = 8'h19;
//assign mul3[8'hff] = 8'h1a;

//assign mul9[8'h00]=8'h00;
//assign mul9[8'h01]=8'h09;
//assign mul9[8'h02]=8'h12;
//assign mul9[8'h03]=8'h1b;
//assign mul9[8'h04]=8'h24;
//assign mul9[8'h05]=8'h2d;
//assign mul9[8'h06]=8'h36;
//assign mul9[8'h07]=8'h3f;
//assign mul9[8'h08]=8'h48;
//assign mul9[8'h09]=8'h41;
//assign mul9[8'h0a]=8'h5a;
//assign mul9[8'h0b]=8'h53;
//assign mul9[8'h0c]=8'h6c;
//assign mul9[8'h0d]=8'h65;
//assign mul9[8'h0e]=8'h7e;
//assign mul9[8'h0f]=8'h77;
//assign mul9[8'h10]=8'h90;
//assign mul9[8'h11]=8'h99;
//assign mul9[8'h12]=8'h82;
//assign mul9[8'h13]=8'h8b;
//assign mul9[8'h14]=8'hb4;
//assign mul9[8'h15]=8'hbd;
//assign mul9[8'h16]=8'ha6;
//assign mul9[8'h17]=8'haf;
//assign mul9[8'h18]=8'hd8;
//assign mul9[8'h19]=8'hd1;
//assign mul9[8'h1a]=8'hca;
//assign mul9[8'h1b]=8'hc3;
//assign mul9[8'h1c]=8'hfc;
//assign mul9[8'h1d]=8'hf5;
//assign mul9[8'h1e]=8'hee;
//assign mul9[8'h1f]=8'he7;
//assign mul9[8'h20]=8'h3b;
//assign mul9[8'h21]=8'h32;
//assign mul9[8'h22]=8'h29;
//assign mul9[8'h23]=8'h20;
//assign mul9[8'h24]=8'h1f;
//assign mul9[8'h25]=8'h16;
//assign mul9[8'h26]=8'h0d;
//assign mul9[8'h27]=8'h04;
//assign mul9[8'h28]=8'h73;
//assign mul9[8'h29]=8'h7a;
//assign mul9[8'h2a]=8'h61;
//assign mul9[8'h2b]=8'h68;
//assign mul9[8'h2c]=8'h57;
//assign mul9[8'h2d]=8'h5e;
//assign mul9[8'h2e]=8'h45;
//assign mul9[8'h2f]=8'h4c;
//assign mul9[8'h30]=8'hab;
//assign mul9[8'h31]=8'ha2;
//assign mul9[8'h32]=8'hb9;
//assign mul9[8'h33]=8'hb0;
//assign mul9[8'h34]=8'h8f;
//assign mul9[8'h35]=8'h86;
//assign mul9[8'h36]=8'h9d;
//assign mul9[8'h37]=8'h94;
//assign mul9[8'h38]=8'he3;
//assign mul9[8'h39]=8'hea;
//assign mul9[8'h3a]=8'hf1;
//assign mul9[8'h3b]=8'hf8;
//assign mul9[8'h3c]=8'hc7;
//assign mul9[8'h3d]=8'hce;
//assign mul9[8'h3e]=8'hd5;
//assign mul9[8'h3f]=8'hdc;
//assign mul9[8'h40]=8'h76;
//assign mul9[8'h41]=8'h7f;
//assign mul9[8'h42]=8'h64;
//assign mul9[8'h43]=8'h6d;
//assign mul9[8'h44]=8'h52;
//assign mul9[8'h45]=8'h5b;
//assign mul9[8'h46]=8'h40;
//assign mul9[8'h47]=8'h49;
//assign mul9[8'h48]=8'h3e;
//assign mul9[8'h49]=8'h37;
//assign mul9[8'h4a]=8'h2c;
//assign mul9[8'h4b]=8'h25;
//assign mul9[8'h4c]=8'h1a;
//assign mul9[8'h4d]=8'h13;
//assign mul9[8'h4e]=8'h08;
//assign mul9[8'h4f]=8'h01;
//assign mul9[8'h50]=8'he6;
//assign mul9[8'h51]=8'hef;
//assign mul9[8'h52]=8'hf4;
//assign mul9[8'h53]=8'hfd;
//assign mul9[8'h54]=8'hc2;
//assign mul9[8'h55]=8'hcb;
//assign mul9[8'h56]=8'hd0;
//assign mul9[8'h57]=8'hd9;
//assign mul9[8'h58]=8'hae;
//assign mul9[8'h59]=8'ha7;
//assign mul9[8'h5a]=8'hbc;
//assign mul9[8'h5b]=8'hb5;
//assign mul9[8'h5c]=8'h8a;
//assign mul9[8'h5d]=8'h83;
//assign mul9[8'h5e]=8'h98;
//assign mul9[8'h5f]=8'h91;
//assign mul9[8'h60]=8'h4d;
//assign mul9[8'h61]=8'h44;
//assign mul9[8'h62]=8'h5f;
//assign mul9[8'h63]=8'h56;
//assign mul9[8'h64]=8'h69;
//assign mul9[8'h65]=8'h60;
//assign mul9[8'h66]=8'h7b;
//assign mul9[8'h67]=8'h72;
//assign mul9[8'h68]=8'h05;
//assign mul9[8'h69]=8'h0c;
//assign mul9[8'h6a]=8'h17;
//assign mul9[8'h6b]=8'h1e;
//assign mul9[8'h6c]=8'h21;
//assign mul9[8'h6d]=8'h28;
//assign mul9[8'h6e]=8'h33;
//assign mul9[8'h6f]=8'h3a;
//assign mul9[8'h70]=8'hdd;
//assign mul9[8'h71]=8'hd4;
//assign mul9[8'h72]=8'hcf;
//assign mul9[8'h73]=8'hc6;
//assign mul9[8'h74]=8'hf9;
//assign mul9[8'h75]=8'hf0;
//assign mul9[8'h76]=8'heb;
//assign mul9[8'h77]=8'he2;
//assign mul9[8'h78]=8'h95;
//assign mul9[8'h79]=8'h9c;
//assign mul9[8'h7a]=8'h87;
//assign mul9[8'h7b]=8'h8e;
//assign mul9[8'h7c]=8'hb1;
//assign mul9[8'h7d]=8'hb8;
//assign mul9[8'h7e]=8'ha3;
//assign mul9[8'h7f]=8'haa;
//assign mul9[8'h80]=8'hec;
//assign mul9[8'h81]=8'he5;
//assign mul9[8'h82]=8'hfe;
//assign mul9[8'h83]=8'hf7;
//assign mul9[8'h84]=8'hc8;
//assign mul9[8'h85]=8'hc1;
//assign mul9[8'h86]=8'hda;
//assign mul9[8'h87]=8'hd3;
//assign mul9[8'h88]=8'ha4;
//assign mul9[8'h89]=8'had;
//assign mul9[8'h8a]=8'hb6;
//assign mul9[8'h8b]=8'hbf;
//assign mul9[8'h8c]=8'h80;
//assign mul9[8'h8d]=8'h89;
//assign mul9[8'h8e]=8'h92;
//assign mul9[8'h8f]=8'h9b;
//assign mul9[8'h90]=8'h7c;
//assign mul9[8'h91]=8'h75;
//assign mul9[8'h92]=8'h6e;
//assign mul9[8'h93]=8'h67;
//assign mul9[8'h94]=8'h58;
//assign mul9[8'h95]=8'h51;
//assign mul9[8'h96]=8'h4a;
//assign mul9[8'h97]=8'h43;
//assign mul9[8'h98]=8'h34;
//assign mul9[8'h99]=8'h3d;
//assign mul9[8'h9a]=8'h26;
//assign mul9[8'h9b]=8'h2f;
//assign mul9[8'h9c]=8'h10;
//assign mul9[8'h9d]=8'h19;
//assign mul9[8'h9e]=8'h02;
//assign mul9[8'h9f]=8'h0b;
//assign mul9[8'ha0]=8'hd7;
//assign mul9[8'ha1]=8'hde;
//assign mul9[8'ha2]=8'hc5;
//assign mul9[8'ha3]=8'hcc;
//assign mul9[8'ha4]=8'hf3;
//assign mul9[8'ha5]=8'hfa;
//assign mul9[8'ha6]=8'he1;
//assign mul9[8'ha7]=8'he8;
//assign mul9[8'ha8]=8'h9f;
//assign mul9[8'ha9]=8'h96;
//assign mul9[8'haa]=8'h8d;
//assign mul9[8'hab]=8'h84;
//assign mul9[8'hac]=8'hbb;
//assign mul9[8'had]=8'hb2;
//assign mul9[8'hae]=8'ha9;
//assign mul9[8'haf]=8'ha0;
//assign mul9[8'hb0]=8'h47;
//assign mul9[8'hb1]=8'h4e;
//assign mul9[8'hb2]=8'h55;
//assign mul9[8'hb3]=8'h5c;
//assign mul9[8'hb4]=8'h63;
//assign mul9[8'hb5]=8'h6a;
//assign mul9[8'hb6]=8'h71;
//assign mul9[8'hb7]=8'h78;
//assign mul9[8'hb8]=8'h0f;
//assign mul9[8'hb9]=8'h06;
//assign mul9[8'hba]=8'h1d;
//assign mul9[8'hbb]=8'h14;
//assign mul9[8'hbc]=8'h2b;
//assign mul9[8'hbd]=8'h22;
//assign mul9[8'hbe]=8'h39;
//assign mul9[8'hbf]=8'h30;
//assign mul9[8'hc0]=8'h9a;
//assign mul9[8'hc1]=8'h93;
//assign mul9[8'hc2]=8'h88;
//assign mul9[8'hc3]=8'h81;
//assign mul9[8'hc4]=8'hbe;
//assign mul9[8'hc5]=8'hb7;
//assign mul9[8'hc6]=8'hac;
//assign mul9[8'hc7]=8'ha5;
//assign mul9[8'hc8]=8'hd2;
//assign mul9[8'hc9]=8'hdb;
//assign mul9[8'hca]=8'hc0;
//assign mul9[8'hcb]=8'hc9;
//assign mul9[8'hcc]=8'hf6;
//assign mul9[8'hcd]=8'hff;
//assign mul9[8'hce]=8'he4;
//assign mul9[8'hcf]=8'hed;
//assign mul9[8'hd0]=8'h0a;
//assign mul9[8'hd1]=8'h03;
//assign mul9[8'hd2]=8'h18;
//assign mul9[8'hd3]=8'h11;
//assign mul9[8'hd4]=8'h2e;
//assign mul9[8'hd5]=8'h27;
//assign mul9[8'hd6]=8'h3c;
//assign mul9[8'hd7]=8'h35;
//assign mul9[8'hd8]=8'h42;
//assign mul9[8'hd9]=8'h4b;
//assign mul9[8'hda]=8'h50;
//assign mul9[8'hdb]=8'h59;
//assign mul9[8'hdc]=8'h66;
//assign mul9[8'hdd]=8'h6f;
//assign mul9[8'hde]=8'h74;
//assign mul9[8'hdf]=8'h7d;
//assign mul9[8'he0]=8'ha1;
//assign mul9[8'he1]=8'ha8;
//assign mul9[8'he2]=8'hb3;
//assign mul9[8'he3]=8'hba;
//assign mul9[8'he4]=8'h85;
//assign mul9[8'he5]=8'h8c;
//assign mul9[8'he6]=8'h97;
//assign mul9[8'he7]=8'h9e;
//assign mul9[8'he8]=8'he9;
//assign mul9[8'he9]=8'he0;
//assign mul9[8'hea]=8'hfb;
//assign mul9[8'heb]=8'hf2;
//assign mul9[8'hec]=8'hcd;
//assign mul9[8'hed]=8'hc4;
//assign mul9[8'hee]=8'hdf;
//assign mul9[8'hef]=8'hd6;
//assign mul9[8'hf0]=8'h31;
//assign mul9[8'hf1]=8'h38;
//assign mul9[8'hf2]=8'h23;
//assign mul9[8'hf3]=8'h2a;
//assign mul9[8'hf4]=8'h15;
//assign mul9[8'hf5]=8'h1c;
//assign mul9[8'hf6]=8'h07;
//assign mul9[8'hf7]=8'h0e;
//assign mul9[8'hf8]=8'h79;
//assign mul9[8'hf9]=8'h70;
//assign mul9[8'hfa]=8'h6b;
//assign mul9[8'hfb]=8'h62;
//assign mul9[8'hfc]=8'h5d;
//assign mul9[8'hfd]=8'h54;
//assign mul9[8'hfe]=8'h4f;
//assign mul9[8'hff]=8'h46;

//assign mul11[8'h00]=8'h00;
//assign mul11[8'h01]=8'h0b;
//assign mul11[8'h02]=8'h16;
//assign mul11[8'h03]=8'h1d;
//assign mul11[8'h04]=8'h2c;
//assign mul11[8'h05]=8'h27;
//assign mul11[8'h06]=8'h3a;
//assign mul11[8'h07]=8'h31;
//assign mul11[8'h08]=8'h58;
//assign mul11[8'h09]=8'h53;
//assign mul11[8'h0a]=8'h4e;
//assign mul11[8'h0b]=8'h45;
//assign mul11[8'h0c]=8'h74;
//assign mul11[8'h0d]=8'h7f;
//assign mul11[8'h0e]=8'h62;
//assign mul11[8'h0f]=8'h69;
//assign mul11[8'h10]=8'hb0;
//assign mul11[8'h11]=8'hbb;
//assign mul11[8'h12]=8'ha6;
//assign mul11[8'h13]=8'had;
//assign mul11[8'h14]=8'h9c;
//assign mul11[8'h15]=8'h97;
//assign mul11[8'h16]=8'h8a;
//assign mul11[8'h17]=8'h81;
//assign mul11[8'h18]=8'he8;
//assign mul11[8'h19]=8'he3;
//assign mul11[8'h1a]=8'hfe;
//assign mul11[8'h1b]=8'hf5;
//assign mul11[8'h1c]=8'hc4;
//assign mul11[8'h1d]=8'hcf;
//assign mul11[8'h1e]=8'hd2;
//assign mul11[8'h1f]=8'hd9;
//assign mul11[8'h20]=8'h7b;
//assign mul11[8'h21]=8'h70;
//assign mul11[8'h22]=8'h6d;
//assign mul11[8'h23]=8'h66;
//assign mul11[8'h24]=8'h57;
//assign mul11[8'h25]=8'h5c;
//assign mul11[8'h26]=8'h41;
//assign mul11[8'h27]=8'h4a;
//assign mul11[8'h28]=8'h23;
//assign mul11[8'h29]=8'h28;
//assign mul11[8'h2a]=8'h35;
//assign mul11[8'h2b]=8'h3e;
//assign mul11[8'h2c]=8'h0f;
//assign mul11[8'h2d]=8'h04;
//assign mul11[8'h2e]=8'h19;
//assign mul11[8'h2f]=8'h12;
//assign mul11[8'h30]=8'hcb;
//assign mul11[8'h31]=8'hc0;
//assign mul11[8'h32]=8'hdd;
//assign mul11[8'h33]=8'hd6;
//assign mul11[8'h34]=8'he7;
//assign mul11[8'h35]=8'hec;
//assign mul11[8'h36]=8'hf1;
//assign mul11[8'h37]=8'hfa;
//assign mul11[8'h38]=8'h93;
//assign mul11[8'h39]=8'h98;
//assign mul11[8'h3a]=8'h85;
//assign mul11[8'h3b]=8'h8e;
//assign mul11[8'h3c]=8'hbf;
//assign mul11[8'h3d]=8'hb4;
//assign mul11[8'h3e]=8'ha9;
//assign mul11[8'h3f]=8'ha2;
//assign mul11[8'h40]=8'hf6;
//assign mul11[8'h41]=8'hfd;
//assign mul11[8'h42]=8'he0;
//assign mul11[8'h43]=8'heb;
//assign mul11[8'h44]=8'hda;
//assign mul11[8'h45]=8'hd1;
//assign mul11[8'h46]=8'hcc;
//assign mul11[8'h47]=8'hc7;
//assign mul11[8'h48]=8'hae;
//assign mul11[8'h49]=8'ha5;
//assign mul11[8'h4a]=8'hb8;
//assign mul11[8'h4b]=8'hb3;
//assign mul11[8'h4c]=8'h82;
//assign mul11[8'h4d]=8'h89;
//assign mul11[8'h4e]=8'h94;
//assign mul11[8'h4f]=8'h9f;
//assign mul11[8'h50]=8'h46;
//assign mul11[8'h51]=8'h4d;
//assign mul11[8'h52]=8'h50;
//assign mul11[8'h53]=8'h5b;
//assign mul11[8'h54]=8'h6a;
//assign mul11[8'h55]=8'h61;
//assign mul11[8'h56]=8'h7c;
//assign mul11[8'h57]=8'h77;
//assign mul11[8'h58]=8'h1e;
//assign mul11[8'h59]=8'h15;
//assign mul11[8'h5a]=8'h08;
//assign mul11[8'h5b]=8'h03;
//assign mul11[8'h5c]=8'h32;
//assign mul11[8'h5d]=8'h39;
//assign mul11[8'h5e]=8'h24;
//assign mul11[8'h5f]=8'h2f;
//assign mul11[8'h60]=8'h8d;
//assign mul11[8'h61]=8'h86;
//assign mul11[8'h62]=8'h9b;
//assign mul11[8'h63]=8'h90;
//assign mul11[8'h64]=8'ha1;
//assign mul11[8'h65]=8'haa;
//assign mul11[8'h66]=8'hb7;
//assign mul11[8'h67]=8'hbc;
//assign mul11[8'h68]=8'hd5;
//assign mul11[8'h69]=8'hde;
//assign mul11[8'h6a]=8'hc3;
//assign mul11[8'h6b]=8'hc8;
//assign mul11[8'h6c]=8'hf9;
//assign mul11[8'h6d]=8'hf2;
//assign mul11[8'h6e]=8'hef;
//assign mul11[8'h6f]=8'he4;
//assign mul11[8'h70]=8'h3d;
//assign mul11[8'h71]=8'h36;
//assign mul11[8'h72]=8'h2b;
//assign mul11[8'h73]=8'h20;
//assign mul11[8'h74]=8'h11;
//assign mul11[8'h75]=8'h1a;
//assign mul11[8'h76]=8'h07;
//assign mul11[8'h77]=8'h0c;
//assign mul11[8'h78]=8'h65;
//assign mul11[8'h79]=8'h6e;
//assign mul11[8'h7a]=8'h73;
//assign mul11[8'h7b]=8'h78;
//assign mul11[8'h7c]=8'h49;
//assign mul11[8'h7d]=8'h42;
//assign mul11[8'h7e]=8'h5f;
//assign mul11[8'h7f]=8'h54;
//assign mul11[8'h80]=8'hf7;
//assign mul11[8'h81]=8'hfc;
//assign mul11[8'h82]=8'he1;
//assign mul11[8'h83]=8'hea;
//assign mul11[8'h84]=8'hdb;
//assign mul11[8'h85]=8'hd0;
//assign mul11[8'h86]=8'hcd;
//assign mul11[8'h87]=8'hc6;
//assign mul11[8'h88]=8'haf;
//assign mul11[8'h89]=8'ha4;
//assign mul11[8'h8a]=8'hb9;
//assign mul11[8'h8b]=8'hb2;
//assign mul11[8'h8c]=8'h83;
//assign mul11[8'h8d]=8'h88;
//assign mul11[8'h8e]=8'h95;
//assign mul11[8'h8f]=8'h9e;
//assign mul11[8'h90]=8'h47;
//assign mul11[8'h91]=8'h4c;
//assign mul11[8'h92]=8'h51;
//assign mul11[8'h93]=8'h5a;
//assign mul11[8'h94]=8'h6b;
//assign mul11[8'h95]=8'h60;
//assign mul11[8'h96]=8'h7d;
//assign mul11[8'h97]=8'h76;
//assign mul11[8'h98]=8'h1f;
//assign mul11[8'h99]=8'h14;
//assign mul11[8'h9a]=8'h09;
//assign mul11[8'h9b]=8'h02;
//assign mul11[8'h9c]=8'h33;
//assign mul11[8'h9d]=8'h38;
//assign mul11[8'h9e]=8'h25;
//assign mul11[8'h9f]=8'h2e;
//assign mul11[8'ha0]=8'h8c;
//assign mul11[8'ha1]=8'h87;
//assign mul11[8'ha2]=8'h9a;
//assign mul11[8'ha3]=8'h91;
//assign mul11[8'ha4]=8'ha0;
//assign mul11[8'ha5]=8'hab;
//assign mul11[8'ha6]=8'hb6;
//assign mul11[8'ha7]=8'hbd;
//assign mul11[8'ha8]=8'hd4;
//assign mul11[8'ha9]=8'hdf;
//assign mul11[8'haa]=8'hc2;
//assign mul11[8'hab]=8'hc9;
//assign mul11[8'hac]=8'hf8;
//assign mul11[8'had]=8'hf3;
//assign mul11[8'hae]=8'hee;
//assign mul11[8'haf]=8'he5;
//assign mul11[8'hb0]=8'h3c;
//assign mul11[8'hb1]=8'h37;
//assign mul11[8'hb2]=8'h2a;
//assign mul11[8'hb3]=8'h21;
//assign mul11[8'hb4]=8'h10;
//assign mul11[8'hb5]=8'h1b;
//assign mul11[8'hb6]=8'h06;
//assign mul11[8'hb7]=8'h0d;
//assign mul11[8'hb8]=8'h64;
//assign mul11[8'hb9]=8'h6f;
//assign mul11[8'hba]=8'h72;
//assign mul11[8'hbb]=8'h79;
//assign mul11[8'hbc]=8'h48;
//assign mul11[8'hbd]=8'h43;
//assign mul11[8'hbe]=8'h5e;
//assign mul11[8'hbf]=8'h55;
//assign mul11[8'hc0]=8'h01;
//assign mul11[8'hc1]=8'h0a;
//assign mul11[8'hc2]=8'h17;
//assign mul11[8'hc3]=8'h1c;
//assign mul11[8'hc4]=8'h2d;
//assign mul11[8'hc5]=8'h26;
//assign mul11[8'hc6]=8'h3b;
//assign mul11[8'hc7]=8'h30;
//assign mul11[8'hc8]=8'h59;
//assign mul11[8'hc9]=8'h52;
//assign mul11[8'hca]=8'h4f;
//assign mul11[8'hcb]=8'h44;
//assign mul11[8'hcc]=8'h75;
//assign mul11[8'hcd]=8'h7e;
//assign mul11[8'hce]=8'h63;
//assign mul11[8'hcf]=8'h68;
//assign mul11[8'hd0]=8'hb1;
//assign mul11[8'hd1]=8'hba;
//assign mul11[8'hd2]=8'ha7;
//assign mul11[8'hd3]=8'hac;
//assign mul11[8'hd4]=8'h9d;
//assign mul11[8'hd5]=8'h96;
//assign mul11[8'hd6]=8'h8b;
//assign mul11[8'hd7]=8'h80;
//assign mul11[8'hd8]=8'he9;
//assign mul11[8'hd9]=8'he2;
//assign mul11[8'hda]=8'hff;
//assign mul11[8'hdb]=8'hf4;
//assign mul11[8'hdc]=8'hc5;
//assign mul11[8'hdd]=8'hce;
//assign mul11[8'hde]=8'hd3;
//assign mul11[8'hdf]=8'hd8;
//assign mul11[8'he0]=8'h7a;
//assign mul11[8'he1]=8'h71;
//assign mul11[8'he2]=8'h6c;
//assign mul11[8'he3]=8'h67;
//assign mul11[8'he4]=8'h56;
//assign mul11[8'he5]=8'h5d;
//assign mul11[8'he6]=8'h40;
//assign mul11[8'he7]=8'h4b;
//assign mul11[8'he8]=8'h22;
//assign mul11[8'he9]=8'h29;
//assign mul11[8'hea]=8'h34;
//assign mul11[8'heb]=8'h3f;
//assign mul11[8'hec]=8'h0e;
//assign mul11[8'hed]=8'h05;
//assign mul11[8'hee]=8'h18;
//assign mul11[8'hef]=8'h13;
//assign mul11[8'hf0]=8'hca;
//assign mul11[8'hf1]=8'hc1;
//assign mul11[8'hf2]=8'hdc;
//assign mul11[8'hf3]=8'hd7;
//assign mul11[8'hf4]=8'he6;
//assign mul11[8'hf5]=8'hed;
//assign mul11[8'hf6]=8'hf0;
//assign mul11[8'hf7]=8'hfb;
//assign mul11[8'hf8]=8'h92;
//assign mul11[8'hf9]=8'h99;
//assign mul11[8'hfa]=8'h84;
//assign mul11[8'hfb]=8'h8f;
//assign mul11[8'hfc]=8'hbe;
//assign mul11[8'hfd]=8'hb5;
//assign mul11[8'hfe]=8'ha8;
//assign mul11[8'hff]=8'ha3;

//assign mul13[8'h00]=8'h00;
//assign mul13[8'h01]=8'h0d;
//assign mul13[8'h02]=8'h1a;
//assign mul13[8'h03]=8'h17;
//assign mul13[8'h04]=8'h34;
//assign mul13[8'h05]=8'h39;
//assign mul13[8'h06]=8'h2e;
//assign mul13[8'h07]=8'h23;
//assign mul13[8'h08]=8'h68;
//assign mul13[8'h09]=8'h65;
//assign mul13[8'h0a]=8'h72;
//assign mul13[8'h0b]=8'h7f;
//assign mul13[8'h0c]=8'h5c;
//assign mul13[8'h0d]=8'h51;
//assign mul13[8'h0e]=8'h46;
//assign mul13[8'h0f]=8'h4b;
//assign mul13[8'h10]=8'hd0;
//assign mul13[8'h11]=8'hdd;
//assign mul13[8'h12]=8'hca;
//assign mul13[8'h13]=8'hc7;
//assign mul13[8'h14]=8'he4;
//assign mul13[8'h15]=8'he9;
//assign mul13[8'h16]=8'hfe;
//assign mul13[8'h17]=8'hf3;
//assign mul13[8'h18]=8'hb8;
//assign mul13[8'h19]=8'hb5;
//assign mul13[8'h1a]=8'ha2;
//assign mul13[8'h1b]=8'haf;
//assign mul13[8'h1c]=8'h8c;
//assign mul13[8'h1d]=8'h81;
//assign mul13[8'h1e]=8'h96;
//assign mul13[8'h1f]=8'h9b;
//assign mul13[8'h20]=8'hbb;
//assign mul13[8'h21]=8'hb6;
//assign mul13[8'h22]=8'ha1;
//assign mul13[8'h23]=8'hac;
//assign mul13[8'h24]=8'h8f;
//assign mul13[8'h25]=8'h82;
//assign mul13[8'h26]=8'h95;
//assign mul13[8'h27]=8'h98;
//assign mul13[8'h28]=8'hd3;
//assign mul13[8'h29]=8'hde;
//assign mul13[8'h2a]=8'hc9;
//assign mul13[8'h2b]=8'hc4;
//assign mul13[8'h2c]=8'he7;
//assign mul13[8'h2d]=8'hea;
//assign mul13[8'h2e]=8'hfd;
//assign mul13[8'h2f]=8'hf0;
//assign mul13[8'h30]=8'h6b;
//assign mul13[8'h31]=8'h66;
//assign mul13[8'h32]=8'h71;
//assign mul13[8'h33]=8'h7c;
//assign mul13[8'h34]=8'h5f;
//assign mul13[8'h35]=8'h52;
//assign mul13[8'h36]=8'h45;
//assign mul13[8'h37]=8'h48;
//assign mul13[8'h38]=8'h03;
//assign mul13[8'h39]=8'h0e;
//assign mul13[8'h3a]=8'h19;
//assign mul13[8'h3b]=8'h14;
//assign mul13[8'h3c]=8'h37;
//assign mul13[8'h3d]=8'h3a;
//assign mul13[8'h3e]=8'h2d;
//assign mul13[8'h3f]=8'h20;
//assign mul13[8'h40]=8'h6d;
//assign mul13[8'h41]=8'h60;
//assign mul13[8'h42]=8'h77;
//assign mul13[8'h43]=8'h7a;
//assign mul13[8'h44]=8'h59;
//assign mul13[8'h45]=8'h54;
//assign mul13[8'h46]=8'h43;
//assign mul13[8'h47]=8'h4e;
//assign mul13[8'h48]=8'h05;
//assign mul13[8'h49]=8'h08;
//assign mul13[8'h4a]=8'h1f;
//assign mul13[8'h4b]=8'h12;
//assign mul13[8'h4c]=8'h31;
//assign mul13[8'h4d]=8'h3c;
//assign mul13[8'h4e]=8'h2b;
//assign mul13[8'h4f]=8'h26;
//assign mul13[8'h50]=8'hbd;
//assign mul13[8'h51]=8'hb0;
//assign mul13[8'h52]=8'ha7;
//assign mul13[8'h53]=8'haa;
//assign mul13[8'h54]=8'h89;
//assign mul13[8'h55]=8'h84;
//assign mul13[8'h56]=8'h93;
//assign mul13[8'h57]=8'h9e;
//assign mul13[8'h58]=8'hd5;
//assign mul13[8'h59]=8'hd8;
//assign mul13[8'h5a]=8'hcf;
//assign mul13[8'h5b]=8'hc2;
//assign mul13[8'h5c]=8'he1;
//assign mul13[8'h5d]=8'hec;
//assign mul13[8'h5e]=8'hfb;
//assign mul13[8'h5f]=8'hf6;
//assign mul13[8'h60]=8'hd6;
//assign mul13[8'h61]=8'hdb;
//assign mul13[8'h62]=8'hcc;
//assign mul13[8'h63]=8'hc1;
//assign mul13[8'h64]=8'he2;
//assign mul13[8'h65]=8'hef;
//assign mul13[8'h66]=8'hf8;
//assign mul13[8'h67]=8'hf5;
//assign mul13[8'h68]=8'hbe;
//assign mul13[8'h69]=8'hb3;
//assign mul13[8'h6a]=8'ha4;
//assign mul13[8'h6b]=8'ha9;
//assign mul13[8'h6c]=8'h8a;
//assign mul13[8'h6d]=8'h87;
//assign mul13[8'h6e]=8'h90;
//assign mul13[8'h6f]=8'h9d;
//assign mul13[8'h70]=8'h06;
//assign mul13[8'h71]=8'h0b;
//assign mul13[8'h72]=8'h1c;
//assign mul13[8'h73]=8'h11;
//assign mul13[8'h74]=8'h32;
//assign mul13[8'h75]=8'h3f;
//assign mul13[8'h76]=8'h28;
//assign mul13[8'h77]=8'h25;
//assign mul13[8'h78]=8'h6e;
//assign mul13[8'h79]=8'h63;
//assign mul13[8'h7a]=8'h74;
//assign mul13[8'h7b]=8'h79;
//assign mul13[8'h7c]=8'h5a;
//assign mul13[8'h7d]=8'h57;
//assign mul13[8'h7e]=8'h40;
//assign mul13[8'h7f]=8'h4d;
//assign mul13[8'h80]=8'hda;
//assign mul13[8'h81]=8'hd7;
//assign mul13[8'h82]=8'hc0;
//assign mul13[8'h83]=8'hcd;
//assign mul13[8'h84]=8'hee;
//assign mul13[8'h85]=8'he3;
//assign mul13[8'h86]=8'hf4;
//assign mul13[8'h87]=8'hf9;
//assign mul13[8'h88]=8'hb2;
//assign mul13[8'h89]=8'hbf;
//assign mul13[8'h8a]=8'ha8;
//assign mul13[8'h8b]=8'ha5;
//assign mul13[8'h8c]=8'h86;
//assign mul13[8'h8d]=8'h8b;
//assign mul13[8'h8e]=8'h9c;
//assign mul13[8'h8f]=8'h91;
//assign mul13[8'h90]=8'h0a;
//assign mul13[8'h91]=8'h07;
//assign mul13[8'h92]=8'h10;
//assign mul13[8'h93]=8'h1d;
//assign mul13[8'h94]=8'h3e;
//assign mul13[8'h95]=8'h33;
//assign mul13[8'h96]=8'h24;
//assign mul13[8'h97]=8'h29;
//assign mul13[8'h98]=8'h62;
//assign mul13[8'h99]=8'h6f;
//assign mul13[8'h9a]=8'h78;
//assign mul13[8'h9b]=8'h75;
//assign mul13[8'h9c]=8'h56;
//assign mul13[8'h9d]=8'h5b;
//assign mul13[8'h9e]=8'h4c;
//assign mul13[8'h9f]=8'h41;
//assign mul13[8'ha0]=8'h61;
//assign mul13[8'ha1]=8'h6c;
//assign mul13[8'ha2]=8'h7b;
//assign mul13[8'ha3]=8'h76;
//assign mul13[8'ha4]=8'h55;
//assign mul13[8'ha5]=8'h58;
//assign mul13[8'ha6]=8'h4f;
//assign mul13[8'ha7]=8'h42;
//assign mul13[8'ha8]=8'h09;
//assign mul13[8'ha9]=8'h04;
//assign mul13[8'haa]=8'h13;
//assign mul13[8'hab]=8'h1e;
//assign mul13[8'hac]=8'h3d;
//assign mul13[8'had]=8'h30;
//assign mul13[8'hae]=8'h27;
//assign mul13[8'haf]=8'h2a;
//assign mul13[8'hb0]=8'hb1;
//assign mul13[8'hb1]=8'hbc;
//assign mul13[8'hb2]=8'hab;
//assign mul13[8'hb3]=8'ha6;
//assign mul13[8'hb4]=8'h85;
//assign mul13[8'hb5]=8'h88;
//assign mul13[8'hb6]=8'h9f;
//assign mul13[8'hb7]=8'h92;
//assign mul13[8'hb8]=8'hd9;
//assign mul13[8'hb9]=8'hd4;
//assign mul13[8'hba]=8'hc3;
//assign mul13[8'hbb]=8'hce;
//assign mul13[8'hbc]=8'hed;
//assign mul13[8'hbd]=8'he0;
//assign mul13[8'hbe]=8'hf7;
//assign mul13[8'hbf]=8'hfa;
//assign mul13[8'hc0]=8'hb7;
//assign mul13[8'hc1]=8'hba;
//assign mul13[8'hc2]=8'had;
//assign mul13[8'hc3]=8'ha0;
//assign mul13[8'hc4]=8'h83;
//assign mul13[8'hc5]=8'h8e;
//assign mul13[8'hc6]=8'h99;
//assign mul13[8'hc7]=8'h94;
//assign mul13[8'hc8]=8'hdf;
//assign mul13[8'hc9]=8'hd2;
//assign mul13[8'hca]=8'hc5;
//assign mul13[8'hcb]=8'hc8;
//assign mul13[8'hcc]=8'heb;
//assign mul13[8'hcd]=8'he6;
//assign mul13[8'hce]=8'hf1;
//assign mul13[8'hcf]=8'hfc;
//assign mul13[8'hd0]=8'h67;
//assign mul13[8'hd1]=8'h6a;
//assign mul13[8'hd2]=8'h7d;
//assign mul13[8'hd3]=8'h70;
//assign mul13[8'hd4]=8'h53;
//assign mul13[8'hd5]=8'h5e;
//assign mul13[8'hd6]=8'h49;
//assign mul13[8'hd7]=8'h44;
//assign mul13[8'hd8]=8'h0f;
//assign mul13[8'hd9]=8'h02;
//assign mul13[8'hda]=8'h15;
//assign mul13[8'hdb]=8'h18;
//assign mul13[8'hdc]=8'h3b;
//assign mul13[8'hdd]=8'h36;
//assign mul13[8'hde]=8'h21;
//assign mul13[8'hdf]=8'h2c;
//assign mul13[8'he0]=8'h0c;
//assign mul13[8'he1]=8'h01;
//assign mul13[8'he2]=8'h16;
//assign mul13[8'he3]=8'h1b;
//assign mul13[8'he4]=8'h38;
//assign mul13[8'he5]=8'h35;
//assign mul13[8'he6]=8'h22;
//assign mul13[8'he7]=8'h2f;
//assign mul13[8'he8]=8'h64;
//assign mul13[8'he9]=8'h69;
//assign mul13[8'hea]=8'h7e;
//assign mul13[8'heb]=8'h73;
//assign mul13[8'hec]=8'h50;
//assign mul13[8'hed]=8'h5d;
//assign mul13[8'hee]=8'h4a;
//assign mul13[8'hef]=8'h47;
//assign mul13[8'hf0]=8'hdc;
//assign mul13[8'hf1]=8'hd1;
//assign mul13[8'hf2]=8'hc6;
//assign mul13[8'hf3]=8'hcb;
//assign mul13[8'hf4]=8'he8;
//assign mul13[8'hf5]=8'he5;
//assign mul13[8'hf6]=8'hf2;
//assign mul13[8'hf7]=8'hff;
//assign mul13[8'hf8]=8'hb4;
//assign mul13[8'hf9]=8'hb9;
//assign mul13[8'hfa]=8'hae;
//assign mul13[8'hfb]=8'ha3;
//assign mul13[8'hfc]=8'h80;
//assign mul13[8'hfd]=8'h8d;
//assign mul13[8'hfe]=8'h9a;
//assign mul13[8'hff]=8'h97;

//assign mul14[8'h00]=8'h00;
//assign mul14[8'h01]=8'h0e;
//assign mul14[8'h02]=8'h1c;
//assign mul14[8'h03]=8'h12;
//assign mul14[8'h04]=8'h38;
//assign mul14[8'h05]=8'h36;
//assign mul14[8'h06]=8'h24;
//assign mul14[8'h07]=8'h2a;
//assign mul14[8'h08]=8'h70;
//assign mul14[8'h09]=8'h7e;
//assign mul14[8'h0a]=8'h6c;
//assign mul14[8'h0b]=8'h62;
//assign mul14[8'h0c]=8'h48;
//assign mul14[8'h0d]=8'h46;
//assign mul14[8'h0e]=8'h54;
//assign mul14[8'h0f]=8'h5a;
//assign mul14[8'h10]=8'he0;
//assign mul14[8'h11]=8'hee;
//assign mul14[8'h12]=8'hfc;
//assign mul14[8'h13]=8'hf2;
//assign mul14[8'h14]=8'hd8;
//assign mul14[8'h15]=8'hd6;
//assign mul14[8'h16]=8'hc4;
//assign mul14[8'h17]=8'hca;
//assign mul14[8'h18]=8'h90;
//assign mul14[8'h19]=8'h9e;
//assign mul14[8'h1a]=8'h8c;
//assign mul14[8'h1b]=8'h82;
//assign mul14[8'h1c]=8'ha8;
//assign mul14[8'h1d]=8'ha6;
//assign mul14[8'h1e]=8'hb4;
//assign mul14[8'h1f]=8'hba;
//assign mul14[8'h20]=8'hdb;
//assign mul14[8'h21]=8'hd5;
//assign mul14[8'h22]=8'hc7;
//assign mul14[8'h23]=8'hc9;
//assign mul14[8'h24]=8'he3;
//assign mul14[8'h25]=8'hed;
//assign mul14[8'h26]=8'hff;
//assign mul14[8'h27]=8'hf1;
//assign mul14[8'h28]=8'hab;
//assign mul14[8'h29]=8'ha5;
//assign mul14[8'h2a]=8'hb7;
//assign mul14[8'h2b]=8'hb9;
//assign mul14[8'h2c]=8'h93;
//assign mul14[8'h2d]=8'h9d;
//assign mul14[8'h2e]=8'h8f;
//assign mul14[8'h2f]=8'h81;
//assign mul14[8'h30]=8'h3b;
//assign mul14[8'h31]=8'h35;
//assign mul14[8'h32]=8'h27;
//assign mul14[8'h33]=8'h29;
//assign mul14[8'h34]=8'h03;
//assign mul14[8'h35]=8'h0d;
//assign mul14[8'h36]=8'h1f;
//assign mul14[8'h37]=8'h11;
//assign mul14[8'h38]=8'h4b;
//assign mul14[8'h39]=8'h45;
//assign mul14[8'h3a]=8'h57;
//assign mul14[8'h3b]=8'h59;
//assign mul14[8'h3c]=8'h73;
//assign mul14[8'h3d]=8'h7d;
//assign mul14[8'h3e]=8'h6f;
//assign mul14[8'h3f]=8'h61;
//assign mul14[8'h40]=8'had;
//assign mul14[8'h41]=8'ha3;
//assign mul14[8'h42]=8'hb1;
//assign mul14[8'h43]=8'hbf;
//assign mul14[8'h44]=8'h95;
//assign mul14[8'h45]=8'h9b;
//assign mul14[8'h46]=8'h89;
//assign mul14[8'h47]=8'h87;
//assign mul14[8'h48]=8'hdd;
//assign mul14[8'h49]=8'hd3;
//assign mul14[8'h4a]=8'hc1;
//assign mul14[8'h4b]=8'hcf;
//assign mul14[8'h4c]=8'he5;
//assign mul14[8'h4d]=8'heb;
//assign mul14[8'h4e]=8'hf9;
//assign mul14[8'h4f]=8'hf7;
//assign mul14[8'h50]=8'h4d;
//assign mul14[8'h51]=8'h43;
//assign mul14[8'h52]=8'h51;
//assign mul14[8'h53]=8'h5f;
//assign mul14[8'h54]=8'h75;
//assign mul14[8'h55]=8'h7b;
//assign mul14[8'h56]=8'h69;
//assign mul14[8'h57]=8'h67;
//assign mul14[8'h58]=8'h3d;
//assign mul14[8'h59]=8'h33;
//assign mul14[8'h5a]=8'h21;
//assign mul14[8'h5b]=8'h2f;
//assign mul14[8'h5c]=8'h05;
//assign mul14[8'h5d]=8'h0b;
//assign mul14[8'h5e]=8'h19;
//assign mul14[8'h5f]=8'h17;
//assign mul14[8'h60]=8'h76;
//assign mul14[8'h61]=8'h78;
//assign mul14[8'h62]=8'h6a;
//assign mul14[8'h63]=8'h64;
//assign mul14[8'h64]=8'h4e;
//assign mul14[8'h65]=8'h40;
//assign mul14[8'h66]=8'h52;
//assign mul14[8'h67]=8'h5c;
//assign mul14[8'h68]=8'h06;
//assign mul14[8'h69]=8'h08;
//assign mul14[8'h6a]=8'h1a;
//assign mul14[8'h6b]=8'h14;
//assign mul14[8'h6c]=8'h3e;
//assign mul14[8'h6d]=8'h30;
//assign mul14[8'h6e]=8'h22;
//assign mul14[8'h6f]=8'h2c;
//assign mul14[8'h70]=8'h96;
//assign mul14[8'h71]=8'h98;
//assign mul14[8'h72]=8'h8a;
//assign mul14[8'h73]=8'h84;
//assign mul14[8'h74]=8'hae;
//assign mul14[8'h75]=8'ha0;
//assign mul14[8'h76]=8'hb2;
//assign mul14[8'h77]=8'hbc;
//assign mul14[8'h78]=8'he6;
//assign mul14[8'h79]=8'he8;
//assign mul14[8'h7a]=8'hfa;
//assign mul14[8'h7b]=8'hf4;
//assign mul14[8'h7c]=8'hde;
//assign mul14[8'h7d]=8'hd0;
//assign mul14[8'h7e]=8'hc2;
//assign mul14[8'h7f]=8'hcc;
//assign mul14[8'h80]=8'h41;
//assign mul14[8'h81]=8'h4f;
//assign mul14[8'h82]=8'h5d;
//assign mul14[8'h83]=8'h53;
//assign mul14[8'h84]=8'h79;
//assign mul14[8'h85]=8'h77;
//assign mul14[8'h86]=8'h65;
//assign mul14[8'h87]=8'h6b;
//assign mul14[8'h88]=8'h31;
//assign mul14[8'h89]=8'h3f;
//assign mul14[8'h8a]=8'h2d;
//assign mul14[8'h8b]=8'h23;
//assign mul14[8'h8c]=8'h09;
//assign mul14[8'h8d]=8'h07;
//assign mul14[8'h8e]=8'h15;
//assign mul14[8'h8f]=8'h1b;
//assign mul14[8'h90]=8'ha1;
//assign mul14[8'h91]=8'haf;
//assign mul14[8'h92]=8'hbd;
//assign mul14[8'h93]=8'hb3;
//assign mul14[8'h94]=8'h99;
//assign mul14[8'h95]=8'h97;
//assign mul14[8'h96]=8'h85;
//assign mul14[8'h97]=8'h8b;
//assign mul14[8'h98]=8'hd1;
//assign mul14[8'h99]=8'hdf;
//assign mul14[8'h9a]=8'hcd;
//assign mul14[8'h9b]=8'hc3;
//assign mul14[8'h9c]=8'he9;
//assign mul14[8'h9d]=8'he7;
//assign mul14[8'h9e]=8'hf5;
//assign mul14[8'h9f]=8'hfb;
//assign mul14[8'ha0]=8'h9a;
//assign mul14[8'ha1]=8'h94;
//assign mul14[8'ha2]=8'h86;
//assign mul14[8'ha3]=8'h88;
//assign mul14[8'ha4]=8'ha2;
//assign mul14[8'ha5]=8'hac;
//assign mul14[8'ha6]=8'hbe;
//assign mul14[8'ha7]=8'hb0;
//assign mul14[8'ha8]=8'hea;
//assign mul14[8'ha9]=8'he4;
//assign mul14[8'haa]=8'hf6;
//assign mul14[8'hab]=8'hf8;
//assign mul14[8'hac]=8'hd2;
//assign mul14[8'had]=8'hdc;
//assign mul14[8'hae]=8'hce;
//assign mul14[8'haf]=8'hc0;
//assign mul14[8'hb0]=8'h7a;
//assign mul14[8'hb1]=8'h74;
//assign mul14[8'hb2]=8'h66;
//assign mul14[8'hb3]=8'h68;
//assign mul14[8'hb4]=8'h42;
//assign mul14[8'hb5]=8'h4c;
//assign mul14[8'hb6]=8'h5e;
//assign mul14[8'hb7]=8'h50;
//assign mul14[8'hb8]=8'h0a;
//assign mul14[8'hb9]=8'h04;
//assign mul14[8'hba]=8'h16;
//assign mul14[8'hbb]=8'h18;
//assign mul14[8'hbc]=8'h32;
//assign mul14[8'hbd]=8'h3c;
//assign mul14[8'hbe]=8'h2e;
//assign mul14[8'hbf]=8'h20;
//assign mul14[8'hc0]=8'hec;
//assign mul14[8'hc1]=8'he2;
//assign mul14[8'hc2]=8'hf0;
//assign mul14[8'hc3]=8'hfe;
//assign mul14[8'hc4]=8'hd4;
//assign mul14[8'hc5]=8'hda;
//assign mul14[8'hc6]=8'hc8;
//assign mul14[8'hc7]=8'hc6;
//assign mul14[8'hc8]=8'h9c;
//assign mul14[8'hc9]=8'h92;
//assign mul14[8'hca]=8'h80;
//assign mul14[8'hcb]=8'h8e;
//assign mul14[8'hcc]=8'ha4;
//assign mul14[8'hcd]=8'haa;
//assign mul14[8'hce]=8'hb8;
//assign mul14[8'hcf]=8'hb6;
//assign mul14[8'hd0]=8'h0c;
//assign mul14[8'hd1]=8'h02;
//assign mul14[8'hd2]=8'h10;
//assign mul14[8'hd3]=8'h1e;
//assign mul14[8'hd4]=8'h34;
//assign mul14[8'hd5]=8'h3a;
//assign mul14[8'hd6]=8'h28;
//assign mul14[8'hd7]=8'h26;
//assign mul14[8'hd8]=8'h7c;
//assign mul14[8'hd9]=8'h72;
//assign mul14[8'hda]=8'h60;
//assign mul14[8'hdb]=8'h6e;
//assign mul14[8'hdc]=8'h44;
//assign mul14[8'hdd]=8'h4a;
//assign mul14[8'hde]=8'h58;
//assign mul14[8'hdf]=8'h56;
//assign mul14[8'he0]=8'h37;
//assign mul14[8'he1]=8'h39;
//assign mul14[8'he2]=8'h2b;
//assign mul14[8'he3]=8'h25;
//assign mul14[8'he4]=8'h0f;
//assign mul14[8'he5]=8'h01;
//assign mul14[8'he6]=8'h13;
//assign mul14[8'he7]=8'h1d;
//assign mul14[8'he8]=8'h47;
//assign mul14[8'he9]=8'h49;
//assign mul14[8'hea]=8'h5b;
//assign mul14[8'heb]=8'h55;
//assign mul14[8'hec]=8'h7f;
//assign mul14[8'hed]=8'h71;
//assign mul14[8'hee]=8'h63;
//assign mul14[8'hef]=8'h6d;
//assign mul14[8'hf0]=8'hd7;
//assign mul14[8'hf1]=8'hd9;
//assign mul14[8'hf2]=8'hcb;
//assign mul14[8'hf3]=8'hc5;
//assign mul14[8'hf4]=8'hef;
//assign mul14[8'hf5]=8'he1;
//assign mul14[8'hf6]=8'hf3;
//assign mul14[8'hf7]=8'hfd;
//assign mul14[8'hf8]=8'ha7;
//assign mul14[8'hf9]=8'ha9;
//assign mul14[8'hfa]=8'hbb;
//assign mul14[8'hfb]=8'hb5;
//assign mul14[8'hfc]=8'h9f;
//assign mul14[8'hfd]=8'h91;
//assign mul14[8'hfe]=8'h83;
//assign mul14[8'hff]=8'h8d;


////assign mcl[127:120]=  (decrypt==0)? ( mul2[a[127:120]] ^ mul3[a[119:112]] ^ a[111:104] ^ a[103:96]):( mul14[a[127:120]] ^ mul11[a[119:112]] ^ mul13[a[111:104]] ^ mul9[a[103:96]]);//state0
////assign mcl[119:112]=  (decrypt==0)? ( a[127:120] ^ mul2[a[119:112]] ^ mul3[a[111:104]] ^ a[103:96]):( mul9[a[127:120]] ^ mul14[a[119:112]] ^ mul11[a[111:104]] ^ mul13[a[103:96]]);//state1
////assign mcl[111:104]=  (decrypt==0)? ( a[127:120] ^ a[119:112] ^ mul2[a[111:104]] ^ mul3[a[103:96]]):( mul13[a[127:120]] ^ mul9[a[119:112]] ^ mul14[a[111:104]] ^ mul11[a[103:96]]);//state2
////assign mcl[103:96]=  (decrypt==0)? ( mul3[a[127:120]] ^ a[119:112] ^ a[111:104] ^ mul2[a[103:96]]):( mul11[a[127:120]] ^ mul13[a[119:112]] ^ mul9[a[111:104]] ^ mul14[a[103:96]]);//state3

////assign mcl[95:88]=   (decrypt==0)? ( mul2[a[95:88]] ^ mul3[a[87:80]] ^ a[79:72] ^ a[71:64]):( mul14[a[95:88]] ^ mul11[a[87:80]] ^ mul13[a[79:72]] ^ mul9[a[71:64]]);//state4
////assign mcl[87:80]=  (decrypt==0)? ( a[95:88] ^ mul2[a[87:80]] ^ mul3[a[79:72]] ^ a[71:64]):( mul9[a[95:88]] ^ mul14[a[87:80]] ^ mul11[a[79:72]] ^ mul13[a[71:64]]);//state5
////assign mcl[79:72]=  (decrypt==0)? ( a[95:88] ^ a[87:80] ^ mul2[a[79:72]] ^ mul3[a[71:64]]):( mul13[a[95:88]] ^ mul9[a[87:80]] ^ mul14[a[79:72]] ^ mul11[a[71:64]]);//state6
////assign mcl[71:64]= (decrypt==0)? ( mul3[a[95:88]] ^ a[87:80] ^ a[79:72] ^ mul2[a[71:64]]):( mul11[a[95:88]] ^ mul13[a[87:80]] ^ mul9[a[79:72]] ^ mul14[a[71:64]]);//state7

////assign mcl[63:56]=  (decrypt==0)? ( mul2[a[63:56]] ^ mul3[a[55:48]] ^ a[47:40] ^ a[39:32]):( mul14[a[63:56]] ^ mul11[a[55:48]] ^ mul13[a[47:40]] ^ mul9[a[39:32]]);//state8
////assign mcl[55:48]=  (decrypt==0)? ( a[63:56] ^ mul2[a[55:48]] ^ mul3[a[47:40]] ^ a[39:32]):( mul9[a[63:56]] ^ mul14[a[55:48]] ^ mul11[a[47:40]] ^ mul13[a[39:32]]);//state9
////assign mcl[47:40]=  (decrypt==0)? ( a[63:56] ^ a[55:48] ^ mul2[a[47:40]] ^ mul3[a[39:32]]):( mul13[a[63:56]] ^ mul9[a[55:48]] ^ mul14[a[47:40]] ^ mul11[a[39:32]]);//state10
////assign mcl[39:32]= (decrypt==0)? ( mul3[a[63:56]] ^ a[55:48] ^ a[47:40] ^ mul2[a[39:32]]):( mul11[a[63:56]] ^ mul13[a[55:48]] ^ mul9[a[47:40]] ^ mul14[a[39:32]]);//state11

////assign mcl[31:24]=  (decrypt==0)? ( mul2[a[31:24]] ^ mul3[a[23:16]] ^ a[15:8] ^ a[7:0]):( mul14[a[31:24]] ^ mul11[a[23:16]] ^ mul13[a[15:8]] ^ mul9[a[7:0]]);//state12
////assign mcl[23:16]=  (decrypt==0)? ( a[31:24] ^ mul2[a[23:16]] ^ mul3[a[15:8]] ^ a[7:0]):( mul9[a[31:24]] ^ mul14[a[23:16]] ^ mul11[a[15:8]] ^ mul13[a[7:0]]);//state13
////assign mcl[15:8]=  (decrypt==0)? ( a[31:24] ^ a[23:16] ^ mul2[a[15:8]] ^ mul3[a[7:0]]):( mul13[a[31:24]] ^ mul9[a[23:16]] ^ mul14[a[15:8]] ^ mul11[a[7:0]]);//state14
////assign mcl[7:0]= (decrypt==0)? ( mul3[a[31:24]] ^ a[23:16] ^ a[15:8] ^ mul2[a[7:0]]):( mul11[a[31:24]] ^ mul13[a[23:16]] ^ mul9[a[15:8]] ^ mul14[a[7:0]]);//state15



//assign mcl[127:120]=  (decrypt==0)? ( mixcolumn32 (a[127:120],a[119:112],a[111:104],a[103:96])):( mul14[a[127:120]] ^ mul11[a[119:112]] ^ mul13[a[111:104]] ^ mul9[a[103:96]]);//state0
//assign mcl[119:112]=  (decrypt==0)? ( mixcolumn32 (a[119:112],a[111:104],a[103:96],a[127:120])):( mul9[a[127:120]] ^ mul14[a[119:112]] ^ mul11[a[111:104]] ^ mul13[a[103:96]]);//state1
//assign mcl[111:104]=  (decrypt==0)? ( mixcolumn32 (a[111:104],a[103:96],a[127:120],a[119:112])):( mul13[a[127:120]] ^ mul9[a[119:112]] ^ mul14[a[111:104]] ^ mul11[a[103:96]]);//state2
//assign mcl[103:96]=  (decrypt==0)? ( mixcolumn32 (a[103:96],a[127:120],a[119:112],a[111:104])):( mul11[a[127:120]] ^ mul13[a[119:112]] ^ mul9[a[111:104]] ^ mul14[a[103:96]]);//state3

//assign mcl[95:88]=   (decrypt==0)? ( mixcolumn32 (a[95:88],a[87:80],a[79:72],a[71:64])):( mul14[a[95:88]] ^ mul11[a[87:80]] ^ mul13[a[79:72]] ^ mul9[a[71:64]]);//state4
//assign mcl[87:80]=  (decrypt==0)? ( mixcolumn32 (a[87:80],a[79:72],a[71:64],a[95:88])):( mul9[a[95:88]] ^ mul14[a[87:80]] ^ mul11[a[79:72]] ^ mul13[a[71:64]]);//state5
//assign mcl[79:72]=  (decrypt==0)? ( mixcolumn32 (a[79:72],a[71:64],a[95:88],a[87:80])):( mul13[a[95:88]] ^ mul9[a[87:80]] ^ mul14[a[79:72]] ^ mul11[a[71:64]]);//state6
//assign mcl[71:64]= (decrypt==0)? ( mixcolumn32 (a[71:64],a[95:88],a[87:80],a[79:72])):( mul11[a[95:88]] ^ mul13[a[87:80]] ^ mul9[a[79:72]] ^ mul14[a[71:64]]);//state7

//assign mcl[63:56]=  (decrypt==0)? ( mixcolumn32 (a[63:56],a[55:48],a[47:40],a[39:32])):( mul14[a[63:56]] ^ mul11[a[55:48]] ^ mul13[a[47:40]] ^ mul9[a[39:32]]);//state8
//assign mcl[55:48]=  (decrypt==0)? ( mixcolumn32 (a[55:48],a[47:40],a[39:32],a[63:56])):( mul9[a[63:56]] ^ mul14[a[55:48]] ^ mul11[a[47:40]] ^ mul13[a[39:32]]);//state9
//assign mcl[47:40]=  (decrypt==0)? ( mixcolumn32 (a[47:40],a[39:32],a[63:56],a[55:48])):( mul13[a[63:56]] ^ mul9[a[55:48]] ^ mul14[a[47:40]] ^ mul11[a[39:32]]);//state10
//assign mcl[39:32]= (decrypt==0)? ( mixcolumn32 (a[39:32],a[63:56],a[55:48],a[47:40])):( mul11[a[63:56]] ^ mul13[a[55:48]] ^ mul9[a[47:40]] ^ mul14[a[39:32]]);//state11

//assign mcl[31:24]=  (decrypt==0)? ( mixcolumn32 (a[31:24],a[23:16],a[15:8],a[7:0])):( mul14[a[31:24]] ^ mul11[a[23:16]] ^ mul13[a[15:8]] ^ mul9[a[7:0]]);//state12
//assign mcl[23:16]=  (decrypt==0)? ( mixcolumn32 (a[23:16],a[15:8],a[7:0],a[31:24])):( mul9[a[31:24]] ^ mul14[a[23:16]] ^ mul11[a[15:8]] ^ mul13[a[7:0]]);//state13
//assign mcl[15:8]=  (decrypt==0)? ( mixcolumn32 (a[15:8],a[7:0],a[31:24],a[23:16])):( mul13[a[31:24]] ^ mul9[a[23:16]] ^ mul14[a[15:8]] ^ mul11[a[7:0]]);//state14
//assign mcl[7:0]= (decrypt==0)? ( mixcolumn32 (a[7:0],a[31:24],a[23:16],a[15:8])):( mul11[a[31:24]] ^ mul13[a[23:16]] ^ mul9[a[15:8]] ^ mul14[a[7:0]]);//state15



////assign mcl[127:120]= mixcolumn32 (a[127:120],a[119:112],a[111:104],a[103:96]);
////assign mcl[119:112]= mixcolumn32 (a[119:112],a[111:104],a[103:96],a[127:120]);
////assign mcl[111:104]= mixcolumn32 (a[111:104],a[103:96],a[127:120],a[119:112]);
////assign mcl[103:96]= mixcolumn32 (a[103:96],a[127:120],a[119:112],a[111:104]);

////assign mcl[95:88]= mixcolumn32 (a[95:88],a[87:80],a[79:72],a[71:64]);
////assign mcl[87:80]= mixcolumn32 (a[87:80],a[79:72],a[71:64],a[95:88]);
////assign mcl[79:72]= mixcolumn32 (a[79:72],a[71:64],a[95:88],a[87:80]);
////assign mcl[71:64]= mixcolumn32 (a[71:64],a[95:88],a[87:80],a[79:72]);

////assign mcl[63:56]= mixcolumn32 (a[63:56],a[55:48],a[47:40],a[39:32]);
////assign mcl[55:48]= mixcolumn32 (a[55:48],a[47:40],a[39:32],a[63:56]);
////assign mcl[47:40]= mixcolumn32 (a[47:40],a[39:32],a[63:56],a[55:48]);
////assign mcl[39:32]= mixcolumn32 (a[39:32],a[63:56],a[55:48],a[47:40]);

////assign mcl[31:24]= mixcolumn32 (a[31:24],a[23:16],a[15:8],a[7:0]);
////assign mcl[23:16]= mixcolumn32 (a[23:16],a[15:8],a[7:0],a[31:24]);
////assign mcl[15:8]= mixcolumn32 (a[15:8],a[7:0],a[31:24],a[23:16]);
////assign mcl[7:0]= mixcolumn32 (a[7:0],a[31:24],a[23:16],a[15:8]);


//function [7:0] mixcolumn32;
//input [7:0] i1,i2,i3,i4;
//begin
//mixcolumn32[7]=i1[6] ^ i2[6] ^ i2[7] ^ i3[7] ^ i4[7];
//mixcolumn32[6]=i1[5] ^ i2[5] ^ i2[6] ^ i3[6] ^ i4[6];
//mixcolumn32[5]=i1[4] ^ i2[4] ^ i2[5] ^ i3[5] ^ i4[5];
//mixcolumn32[4]=i1[3] ^ i1[7] ^ i2[3] ^ i2[4] ^ i2[7] ^ i3[4] ^ i4[4];
//mixcolumn32[3]=i1[2] ^ i1[7] ^ i2[2] ^ i2[3] ^ i2[7] ^ i3[3] ^ i4[3];
//mixcolumn32[2]=i1[1] ^ i2[1] ^ i2[2] ^ i3[2] ^ i4[2];
//mixcolumn32[1]=i1[0] ^ i1[7] ^ i2[0] ^ i2[1] ^ i2[7] ^ i3[1] ^ i4[1];
//mixcolumn32[0]=i1[7] ^ i2[7] ^ i2[0] ^ i3[0] ^ i4[0];
//end
//endfunction


//----------------------------------------------------------------
// Gaolis multiplication functions for Inverse MixColumn.
//----------------------------------------------------------------
function [7 : 0] gm2(input [7 : 0] op);
begin
  gm2 = {op[6 : 0], 1'b0} ^ (8'h1b & {8{op[7]}});
end
endfunction // gm2

function [7 : 0] gm3(input [7 : 0] op);
begin
  gm3 = gm2(op) ^ op;
end
endfunction // gm3

function [7 : 0] gm4(input [7 : 0] op);
begin
  gm4 = gm2(gm2(op));
end
endfunction // gm4

function [7 : 0] gm8(input [7 : 0] op);
begin
  gm8 = gm2(gm4(op));
end
endfunction // gm8

function [7 : 0] gm09(input [7 : 0] op);
begin
  gm09 = gm8(op) ^ op;
end
endfunction // gm09

function [7 : 0] gm11(input [7 : 0] op);
begin
  gm11 = gm8(op) ^ gm2(op) ^ op;
end
endfunction // gm11

function [7 : 0] gm13(input [7 : 0] op);
begin
  gm13 = gm8(op) ^ gm4(op) ^ op;
end
endfunction // gm13

function [7 : 0] gm14(input [7 : 0] op);
begin
  gm14 = gm8(op) ^ gm4(op) ^ gm2(op);
end
endfunction // gm14

function [31 : 0] inv_mixw(input [31 : 0] w);
reg [7 : 0] b0, b1, b2, b3;
reg [7 : 0] mb0, mb1, mb2, mb3;
begin
  b0 = w[31 : 24];
  b1 = w[23 : 16];
  b2 = w[15 : 08];
  b3 = w[07 : 00];

  mb0 = gm14(b0) ^ gm11(b1) ^ gm13(b2) ^ gm09(b3);
  mb1 = gm09(b0) ^ gm14(b1) ^ gm11(b2) ^ gm13(b3);
  mb2 = gm13(b0) ^ gm09(b1) ^ gm14(b2) ^ gm11(b3);
  mb3 = gm11(b0) ^ gm13(b1) ^ gm09(b2) ^ gm14(b3);

  inv_mixw = {mb0, mb1, mb2, mb3};
end
endfunction // mixw

function [127 : 0] inv_mixcolumns(input [127 : 0] data);
reg [31 : 0] w0, w1, w2, w3;
reg [31 : 0] ws0, ws1, ws2, ws3;
begin
  w0 = data[127 : 096];
  w1 = data[095 : 064];
  w2 = data[063 : 032];
  w3 = data[031 : 000];

  ws0 = inv_mixw(w0);
  ws1 = inv_mixw(w1);
  ws2 = inv_mixw(w2);
  ws3 = inv_mixw(w3);

  inv_mixcolumns = {ws0, ws1, ws2, ws3};
end
endfunction // inv_mixcolumns


function [31 : 0] mixw(input [31 : 0] w);
reg [7 : 0] b0, b1, b2, b3;
reg [7 : 0] mb0, mb1, mb2, mb3;
begin
  b0 = w[31 : 24];
  b1 = w[23 : 16];
  b2 = w[15 : 08];
  b3 = w[07 : 00];

  mb0 = gm2(b0) ^ gm3(b1) ^ b2      ^ b3;
  mb1 = b0      ^ gm2(b1) ^ gm3(b2) ^ b3;
  mb2 = b0      ^ b1      ^ gm2(b2) ^ gm3(b3);
  mb3 = gm3(b0) ^ b1      ^ b2      ^ gm2(b3);

  mixw = {mb0, mb1, mb2, mb3};
end
endfunction // mixw

function [127 : 0] mixcolumns(input [127 : 0] data);
reg [31 : 0] w0, w1, w2, w3;
reg [31 : 0] ws0, ws1, ws2, ws3;
begin
  w0 = data[127 : 096];
  w1 = data[095 : 064];
  w2 = data[063 : 032];
  w3 = data[031 : 000];

  ws0 = mixw(w0);
  ws1 = mixw(w1);
  ws2 = mixw(w2);
  ws3 = mixw(w3);

  mixcolumns = {ws0, ws1, ws2, ws3};
end
endfunction // mixcolumns



endmodule
